parameter sim_test = "random" ; 
        parameter nums = 30;
        parameter max_delay = 5;  // run test
