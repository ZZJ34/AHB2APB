task display_name();
  $display("Starting    %s task !!!", name);
endtask

task transfer_AHB_trans(input nums=0);
    i_apb_if.haddr = {`HADDR_SYS_WIDTH{1'b1}};
endtask
